`ifdef VERILATOR
	`define SIMULATION   // for verilator simulation only
`endif

module Tx_top
(clk, 
`ifdef SIMULATION
	start, i_data,
`endif
serial_out);   // UART transmitter :  parallel input, serial output (PISO)

input clk;  // 48MHz
// input reset;  // will be added later to clear various registers

`ifdef SIMULATION
	input start;     // i_data is valid, so start transmission. This 'start' signal is set to '1' for one baud clock cycle
	input[7:0] i_data; 	// parallel input
`else
	wire[7:0] i_data = 8'h46; 	// equivalent ASCII code in hex radix for the character 'F'
`endif

output serial_out;  // serial output from serializer (TxUART)

wire baud_clk;  // 9600bps baudrate clock
wire enable;   	// starts transmission or not
wire o_busy, start_tx, parity_bit;

TxUART tx (.clk(clk), .baud_clk(baud_clk), .enable(enable), .i_data(i_data), .o_busy(o_busy), .start_tx(start_tx));

baud_generator bg (.clk(clk), .baud_clk(baud_clk));	// to derive the desired baud rate of 9600bps

`ifdef SIMULATION
	assign enable = start;
`else
	enable_generator eg (.clk(clk), .en_out(enable));   // transmission is enabled/repeated every 500ms
`endif
	
shift_register PISO (.clk(baud_clk), .valid(start_tx), .tx_busy(o_busy), .data_in({parity_bit, i_data}), .data_out(serial_out)); // .data_in({parity_bit, i_data  --> transmit LSB first

// FIFO tx_fifo (clk, reset, enqueue, dequeue, flush, i_value, almost_full, almost_empty, o_value);

assign parity_bit = ^i_data; // even parity http://www.asic-world.com/examples/verilog/parity.html

endmodule
