module shift_register(clk, valid, tx_busy, data_in, data_out);   // PISO shift register specificaly for UART Tx

input clk, valid, tx_busy;	// clock, data is valid, tx is not in idle state
input [8:0] data_in;   // parallel input, 8-bits data + 1-bit parity
output reg data_out;	// serial output

reg [8:0] data_shift_reg;
//integer index=0;
always @(posedge clk)
begin
    if (valid && (!tx_busy))   // only accept input data when Tx is in idle state and data is valid	 
	data_shift_reg <= data_in;   // prepare to start shifting in new chunk of data
    else
	data_shift_reg <= { 1'b1, data_shift_reg[8:1] };   // pushes 1 in such that when tx finishes, a logic level of '1' is transmitted
end

always @(posedge clk)
begin
    if (valid && (!tx_busy)) begin	// only start shifting out data when Tx is in idle state and data is valid
	data_out <= 1'b0;  // 0-bit represents UART start bit
	//$display("UART start bit = %1b, time = %f", data_out, $realtime);
    end
    else if (tx_busy) begin
	data_out <= data_shift_reg[0];  // transmit LSB first according to UART protocol
	//$display("UART data bit[%1d] = %1b, time = %f", index, data_out, $realtime); index = index + 1;
    end
    else
	data_out <= 1'b1;  // UART Tx line is pulled HIGH as default to signal IDLING state both *before* and *after* UART transmission
end

endmodule
